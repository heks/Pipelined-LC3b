--
-- VHDL Architecture ece411.ZEXTLowerB1.untitled
--
-- Created:
--          by - labelle1.ews (siebl-0220-08.ews.illinois.edu)
--          at - 00:28:53 04/12/13
--
-- using Mentor Graphics HDL Designer(TM) 2012.1 (Build 6)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.NUMERIC_STD.all;

LIBRARY ece411;
USE ece411.LC3b_types.all;

ENTITY ZEXTLowerB1 IS
-- Declarations

END ZEXTLowerB1 ;

--
ARCHITECTURE untitled OF ZEXTLowerB1 IS
BEGIN
END ARCHITECTURE untitled;

